../../../scramble_rel001_papilio/source/scramble_dblscan.vhd