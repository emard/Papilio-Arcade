../../../scramble_rel001_papilio/source/T80/T80_Reg.vhd